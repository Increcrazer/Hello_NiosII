// hello.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module hello (
		input  wire  clk_0_clk,     // clk_0.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] cpu_0_data_master_readdata;                                // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_waitrequest;                             // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire         cpu_0_data_master_debugaccess;                             // cpu_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire  [18:0] cpu_0_data_master_address;                                 // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;                              // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_0_data_master_read;                                    // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire         cpu_0_data_master_write;                                   // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                               // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [31:0] cpu_0_instruction_master_readdata;                         // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;                      // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [18:0] cpu_0_instruction_master_address;                          // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                             // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_readdata;        // cpu_0:jtag_debug_module_readdata -> mm_interconnect_0:cpu_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest;     // cpu_0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess;     // mm_interconnect_0:cpu_0_jtag_debug_module_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_0_jtag_debug_module_address;         // mm_interconnect_0:cpu_0_jtag_debug_module_address -> cpu_0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_read;            // mm_interconnect_0:cpu_0_jtag_debug_module_read -> cpu_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_0_jtag_debug_module_byteenable;      // mm_interconnect_0:cpu_0_jtag_debug_module_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_write;           // mm_interconnect_0:cpu_0_jtag_debug_module_write -> cpu_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_writedata;       // mm_interconnect_0:cpu_0_jtag_debug_module_writedata -> cpu_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_0_d_irq_irq;                                           // irq_mapper:sender_irq -> cpu_0:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu_0:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_0_reset_n_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [onchip_memory2:reset_req, rst_translator_001:reset_req_in]
	wire         cpu_0_jtag_debug_module_reset_reset;                       // cpu_0:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1

	hello_cpu_0 cpu_0 (
		.clk                                   (clk_0_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (cpu_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                               //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	hello_jtag_uart jtag_uart (
		.clk            (clk_0_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	hello_onchip_memory2 onchip_memory2 (
		.clk        (clk_0_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	hello_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_0_clk),                                                 //                             clk_0_clk.clk
		.cpu_0_reset_n_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            //   cpu_0_reset_n_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // jtag_uart_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                   (cpu_0_data_master_address),                                 //                     cpu_0_data_master.address
		.cpu_0_data_master_waitrequest               (cpu_0_data_master_waitrequest),                             //                                      .waitrequest
		.cpu_0_data_master_byteenable                (cpu_0_data_master_byteenable),                              //                                      .byteenable
		.cpu_0_data_master_read                      (cpu_0_data_master_read),                                    //                                      .read
		.cpu_0_data_master_readdata                  (cpu_0_data_master_readdata),                                //                                      .readdata
		.cpu_0_data_master_write                     (cpu_0_data_master_write),                                   //                                      .write
		.cpu_0_data_master_writedata                 (cpu_0_data_master_writedata),                               //                                      .writedata
		.cpu_0_data_master_debugaccess               (cpu_0_data_master_debugaccess),                             //                                      .debugaccess
		.cpu_0_instruction_master_address            (cpu_0_instruction_master_address),                          //              cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest        (cpu_0_instruction_master_waitrequest),                      //                                      .waitrequest
		.cpu_0_instruction_master_read               (cpu_0_instruction_master_read),                             //                                      .read
		.cpu_0_instruction_master_readdata           (cpu_0_instruction_master_readdata),                         //                                      .readdata
		.cpu_0_jtag_debug_module_address             (mm_interconnect_0_cpu_0_jtag_debug_module_address),         //               cpu_0_jtag_debug_module.address
		.cpu_0_jtag_debug_module_write               (mm_interconnect_0_cpu_0_jtag_debug_module_write),           //                                      .write
		.cpu_0_jtag_debug_module_read                (mm_interconnect_0_cpu_0_jtag_debug_module_read),            //                                      .read
		.cpu_0_jtag_debug_module_readdata            (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),        //                                      .readdata
		.cpu_0_jtag_debug_module_writedata           (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),       //                                      .writedata
		.cpu_0_jtag_debug_module_byteenable          (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),      //                                      .byteenable
		.cpu_0_jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest),     //                                      .waitrequest
		.cpu_0_jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess),     //                                      .debugaccess
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.onchip_memory2_s1_address                   (mm_interconnect_0_onchip_memory2_s1_address),               //                     onchip_memory2_s1.address
		.onchip_memory2_s1_write                     (mm_interconnect_0_onchip_memory2_s1_write),                 //                                      .write
		.onchip_memory2_s1_readdata                  (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                      .readdata
		.onchip_memory2_s1_writedata                 (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                      .writedata
		.onchip_memory2_s1_byteenable                (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                      .byteenable
		.onchip_memory2_s1_chipselect                (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                      .chipselect
		.onchip_memory2_s1_clken                     (mm_interconnect_0_onchip_memory2_s1_clken)                  //                                      .clken
	);

	hello_irq_mapper irq_mapper (
		.clk           (clk_0_clk),                      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_0_clk),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_0_jtag_debug_module_reset_reset),    // reset_in1.reset
		.clk            (clk_0_clk),                              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
