
module hello (
	clk_0_clk,
	reset_reset_n);	

	input		clk_0_clk;
	input		reset_reset_n;
endmodule
